// nios_led3.v

// Generated using ACDS version 23.1 991

`timescale 1 ps / 1 ps
module nios_led3 (
		input  wire        clk_clk,         //      clk.clk
		input  wire [1:0]  i_btn_export,    //    i_btn.export
		input  wire [9:0]  i_switch_export, // i_switch.export
		output wire [1:0]  o_ledr_export,   //   o_ledr.export
		output wire [31:0] o_sseg_export,   //   o_sseg.export
		input  wire        reset_reset_n    //    reset.reset_n
	);

	wire  [31:0] cpu_nios_led3_data_master_readdata;                          // mm_interconnect_0:cpu_nios_led3_data_master_readdata -> cpu_nios_led3:d_readdata
	wire         cpu_nios_led3_data_master_waitrequest;                       // mm_interconnect_0:cpu_nios_led3_data_master_waitrequest -> cpu_nios_led3:d_waitrequest
	wire         cpu_nios_led3_data_master_debugaccess;                       // cpu_nios_led3:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:cpu_nios_led3_data_master_debugaccess
	wire  [18:0] cpu_nios_led3_data_master_address;                           // cpu_nios_led3:d_address -> mm_interconnect_0:cpu_nios_led3_data_master_address
	wire   [3:0] cpu_nios_led3_data_master_byteenable;                        // cpu_nios_led3:d_byteenable -> mm_interconnect_0:cpu_nios_led3_data_master_byteenable
	wire         cpu_nios_led3_data_master_read;                              // cpu_nios_led3:d_read -> mm_interconnect_0:cpu_nios_led3_data_master_read
	wire         cpu_nios_led3_data_master_write;                             // cpu_nios_led3:d_write -> mm_interconnect_0:cpu_nios_led3_data_master_write
	wire  [31:0] cpu_nios_led3_data_master_writedata;                         // cpu_nios_led3:d_writedata -> mm_interconnect_0:cpu_nios_led3_data_master_writedata
	wire  [31:0] cpu_nios_led3_instruction_master_readdata;                   // mm_interconnect_0:cpu_nios_led3_instruction_master_readdata -> cpu_nios_led3:i_readdata
	wire         cpu_nios_led3_instruction_master_waitrequest;                // mm_interconnect_0:cpu_nios_led3_instruction_master_waitrequest -> cpu_nios_led3:i_waitrequest
	wire  [18:0] cpu_nios_led3_instruction_master_address;                    // cpu_nios_led3:i_address -> mm_interconnect_0:cpu_nios_led3_instruction_master_address
	wire         cpu_nios_led3_instruction_master_read;                       // cpu_nios_led3:i_read -> mm_interconnect_0:cpu_nios_led3_instruction_master_read
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;    // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;      // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest;   // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;       // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;          // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;         // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;     // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire  [31:0] mm_interconnect_0_cpu_nios_led3_debug_mem_slave_readdata;    // cpu_nios_led3:debug_mem_slave_readdata -> mm_interconnect_0:cpu_nios_led3_debug_mem_slave_readdata
	wire         mm_interconnect_0_cpu_nios_led3_debug_mem_slave_waitrequest; // cpu_nios_led3:debug_mem_slave_waitrequest -> mm_interconnect_0:cpu_nios_led3_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_cpu_nios_led3_debug_mem_slave_debugaccess; // mm_interconnect_0:cpu_nios_led3_debug_mem_slave_debugaccess -> cpu_nios_led3:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_cpu_nios_led3_debug_mem_slave_address;     // mm_interconnect_0:cpu_nios_led3_debug_mem_slave_address -> cpu_nios_led3:debug_mem_slave_address
	wire         mm_interconnect_0_cpu_nios_led3_debug_mem_slave_read;        // mm_interconnect_0:cpu_nios_led3_debug_mem_slave_read -> cpu_nios_led3:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_cpu_nios_led3_debug_mem_slave_byteenable;  // mm_interconnect_0:cpu_nios_led3_debug_mem_slave_byteenable -> cpu_nios_led3:debug_mem_slave_byteenable
	wire         mm_interconnect_0_cpu_nios_led3_debug_mem_slave_write;       // mm_interconnect_0:cpu_nios_led3_debug_mem_slave_write -> cpu_nios_led3:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_cpu_nios_led3_debug_mem_slave_writedata;   // mm_interconnect_0:cpu_nios_led3_debug_mem_slave_writedata -> cpu_nios_led3:debug_mem_slave_writedata
	wire         mm_interconnect_0_ram_s1_chipselect;                         // mm_interconnect_0:RAM_s1_chipselect -> RAM:chipselect
	wire  [31:0] mm_interconnect_0_ram_s1_readdata;                           // RAM:readdata -> mm_interconnect_0:RAM_s1_readdata
	wire  [14:0] mm_interconnect_0_ram_s1_address;                            // mm_interconnect_0:RAM_s1_address -> RAM:address
	wire   [3:0] mm_interconnect_0_ram_s1_byteenable;                         // mm_interconnect_0:RAM_s1_byteenable -> RAM:byteenable
	wire         mm_interconnect_0_ram_s1_write;                              // mm_interconnect_0:RAM_s1_write -> RAM:write
	wire  [31:0] mm_interconnect_0_ram_s1_writedata;                          // mm_interconnect_0:RAM_s1_writedata -> RAM:writedata
	wire         mm_interconnect_0_ram_s1_clken;                              // mm_interconnect_0:RAM_s1_clken -> RAM:clken
	wire  [31:0] mm_interconnect_0_switch_s1_readdata;                        // switch:readdata -> mm_interconnect_0:switch_s1_readdata
	wire   [1:0] mm_interconnect_0_switch_s1_address;                         // mm_interconnect_0:switch_s1_address -> switch:address
	wire         mm_interconnect_0_btn_s1_chipselect;                         // mm_interconnect_0:btn_s1_chipselect -> btn:chipselect
	wire  [31:0] mm_interconnect_0_btn_s1_readdata;                           // btn:readdata -> mm_interconnect_0:btn_s1_readdata
	wire   [1:0] mm_interconnect_0_btn_s1_address;                            // mm_interconnect_0:btn_s1_address -> btn:address
	wire         mm_interconnect_0_btn_s1_write;                              // mm_interconnect_0:btn_s1_write -> btn:write_n
	wire  [31:0] mm_interconnect_0_btn_s1_writedata;                          // mm_interconnect_0:btn_s1_writedata -> btn:writedata
	wire         mm_interconnect_0_ledr_s1_chipselect;                        // mm_interconnect_0:ledr_s1_chipselect -> ledr:chipselect
	wire  [31:0] mm_interconnect_0_ledr_s1_readdata;                          // ledr:readdata -> mm_interconnect_0:ledr_s1_readdata
	wire   [1:0] mm_interconnect_0_ledr_s1_address;                           // mm_interconnect_0:ledr_s1_address -> ledr:address
	wire         mm_interconnect_0_ledr_s1_write;                             // mm_interconnect_0:ledr_s1_write -> ledr:write_n
	wire  [31:0] mm_interconnect_0_ledr_s1_writedata;                         // mm_interconnect_0:ledr_s1_writedata -> ledr:writedata
	wire         mm_interconnect_0_sseg_s1_chipselect;                        // mm_interconnect_0:sseg_s1_chipselect -> sseg:chipselect
	wire  [31:0] mm_interconnect_0_sseg_s1_readdata;                          // sseg:readdata -> mm_interconnect_0:sseg_s1_readdata
	wire   [1:0] mm_interconnect_0_sseg_s1_address;                           // mm_interconnect_0:sseg_s1_address -> sseg:address
	wire         mm_interconnect_0_sseg_s1_write;                             // mm_interconnect_0:sseg_s1_write -> sseg:write_n
	wire  [31:0] mm_interconnect_0_sseg_s1_writedata;                         // mm_interconnect_0:sseg_s1_writedata -> sseg:writedata
	wire         mm_interconnect_0_sys_timer_s1_chipselect;                   // mm_interconnect_0:sys_timer_s1_chipselect -> sys_timer:chipselect
	wire  [15:0] mm_interconnect_0_sys_timer_s1_readdata;                     // sys_timer:readdata -> mm_interconnect_0:sys_timer_s1_readdata
	wire   [2:0] mm_interconnect_0_sys_timer_s1_address;                      // mm_interconnect_0:sys_timer_s1_address -> sys_timer:address
	wire         mm_interconnect_0_sys_timer_s1_write;                        // mm_interconnect_0:sys_timer_s1_write -> sys_timer:write_n
	wire  [15:0] mm_interconnect_0_sys_timer_s1_writedata;                    // mm_interconnect_0:sys_timer_s1_writedata -> sys_timer:writedata
	wire         mm_interconnect_0_usr_timer_s1_chipselect;                   // mm_interconnect_0:usr_timer_s1_chipselect -> usr_timer:chipselect
	wire  [15:0] mm_interconnect_0_usr_timer_s1_readdata;                     // usr_timer:readdata -> mm_interconnect_0:usr_timer_s1_readdata
	wire   [2:0] mm_interconnect_0_usr_timer_s1_address;                      // mm_interconnect_0:usr_timer_s1_address -> usr_timer:address
	wire         mm_interconnect_0_usr_timer_s1_write;                        // mm_interconnect_0:usr_timer_s1_write -> usr_timer:write_n
	wire  [15:0] mm_interconnect_0_usr_timer_s1_writedata;                    // mm_interconnect_0:usr_timer_s1_writedata -> usr_timer:writedata
	wire         irq_mapper_receiver0_irq;                                    // btn:irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                    // sys_timer:irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                    // usr_timer:irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                                    // jtag_uart:av_irq -> irq_mapper:receiver3_irq
	wire  [31:0] cpu_nios_led3_irq_irq;                                       // irq_mapper:sender_irq -> cpu_nios_led3:irq
	wire         rst_controller_reset_out_reset;                              // rst_controller:reset_out -> [RAM:reset, btn:reset_n, cpu_nios_led3:reset_n, irq_mapper:reset, jtag_uart:rst_n, ledr:reset_n, mm_interconnect_0:cpu_nios_led3_reset_reset_bridge_in_reset_reset, rst_translator:in_reset, sseg:reset_n, switch:reset_n, sys_timer:reset_n, usr_timer:reset_n]
	wire         rst_controller_reset_out_reset_req;                          // rst_controller:reset_req -> [RAM:reset_req, cpu_nios_led3:reset_req, rst_translator:reset_req_in]

	nios_led3_RAM ram (
		.clk        (clk_clk),                             //   clk1.clk
		.address    (mm_interconnect_0_ram_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_ram_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_ram_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_ram_s1_write),      //       .write
		.readdata   (mm_interconnect_0_ram_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_ram_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_ram_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),      // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),  //       .reset_req
		.freeze     (1'b0)                                 // (terminated)
	);

	nios_led3_btn btn (
		.clk        (clk_clk),                             //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_0_btn_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_btn_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_btn_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_btn_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_btn_s1_readdata),   //                    .readdata
		.in_port    (i_btn_export),                        // external_connection.export
		.irq        (irq_mapper_receiver0_irq)             //                 irq.irq
	);

	nios_led3_cpu_nios_led3 cpu_nios_led3 (
		.clk                                 (clk_clk),                                                     //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                             //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                          //                          .reset_req
		.d_address                           (cpu_nios_led3_data_master_address),                           //               data_master.address
		.d_byteenable                        (cpu_nios_led3_data_master_byteenable),                        //                          .byteenable
		.d_read                              (cpu_nios_led3_data_master_read),                              //                          .read
		.d_readdata                          (cpu_nios_led3_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (cpu_nios_led3_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (cpu_nios_led3_data_master_write),                             //                          .write
		.d_writedata                         (cpu_nios_led3_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (cpu_nios_led3_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (cpu_nios_led3_instruction_master_address),                    //        instruction_master.address
		.i_read                              (cpu_nios_led3_instruction_master_read),                       //                          .read
		.i_readdata                          (cpu_nios_led3_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (cpu_nios_led3_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (cpu_nios_led3_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (),                                                            //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_cpu_nios_led3_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_cpu_nios_led3_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_cpu_nios_led3_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_cpu_nios_led3_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_cpu_nios_led3_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_cpu_nios_led3_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_cpu_nios_led3_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_cpu_nios_led3_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                             // custom_instruction_master.readra
	);

	nios_led3_jtag_uart jtag_uart (
		.clk            (clk_clk),                                                   //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                           //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver3_irq)                                   //               irq.irq
	);

	nios_led3_ledr ledr (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_ledr_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_ledr_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_ledr_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_ledr_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_ledr_s1_readdata),   //                    .readdata
		.out_port   (o_ledr_export)                         // external_connection.export
	);

	nios_led3_sseg sseg (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_sseg_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_sseg_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_sseg_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_sseg_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_sseg_s1_readdata),   //                    .readdata
		.out_port   (o_sseg_export)                         // external_connection.export
	);

	nios_led3_switch switch (
		.clk      (clk_clk),                              //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address  (mm_interconnect_0_switch_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_switch_s1_readdata), //                    .readdata
		.in_port  (i_switch_export)                       // external_connection.export
	);

	nios_led3_sys_timer sys_timer (
		.clk        (clk_clk),                                   //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           // reset.reset_n
		.address    (mm_interconnect_0_sys_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_sys_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_sys_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_sys_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_sys_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver1_irq)                   //   irq.irq
	);

	nios_led3_sys_timer usr_timer (
		.clk        (clk_clk),                                   //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           // reset.reset_n
		.address    (mm_interconnect_0_usr_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_usr_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_usr_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_usr_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_usr_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver2_irq)                   //   irq.irq
	);

	nios_led3_mm_interconnect_0 mm_interconnect_0 (
		.clk_clk_clk                                     (clk_clk),                                                     //                                   clk_clk.clk
		.cpu_nios_led3_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                              // cpu_nios_led3_reset_reset_bridge_in_reset.reset
		.cpu_nios_led3_data_master_address               (cpu_nios_led3_data_master_address),                           //                 cpu_nios_led3_data_master.address
		.cpu_nios_led3_data_master_waitrequest           (cpu_nios_led3_data_master_waitrequest),                       //                                          .waitrequest
		.cpu_nios_led3_data_master_byteenable            (cpu_nios_led3_data_master_byteenable),                        //                                          .byteenable
		.cpu_nios_led3_data_master_read                  (cpu_nios_led3_data_master_read),                              //                                          .read
		.cpu_nios_led3_data_master_readdata              (cpu_nios_led3_data_master_readdata),                          //                                          .readdata
		.cpu_nios_led3_data_master_write                 (cpu_nios_led3_data_master_write),                             //                                          .write
		.cpu_nios_led3_data_master_writedata             (cpu_nios_led3_data_master_writedata),                         //                                          .writedata
		.cpu_nios_led3_data_master_debugaccess           (cpu_nios_led3_data_master_debugaccess),                       //                                          .debugaccess
		.cpu_nios_led3_instruction_master_address        (cpu_nios_led3_instruction_master_address),                    //          cpu_nios_led3_instruction_master.address
		.cpu_nios_led3_instruction_master_waitrequest    (cpu_nios_led3_instruction_master_waitrequest),                //                                          .waitrequest
		.cpu_nios_led3_instruction_master_read           (cpu_nios_led3_instruction_master_read),                       //                                          .read
		.cpu_nios_led3_instruction_master_readdata       (cpu_nios_led3_instruction_master_readdata),                   //                                          .readdata
		.btn_s1_address                                  (mm_interconnect_0_btn_s1_address),                            //                                    btn_s1.address
		.btn_s1_write                                    (mm_interconnect_0_btn_s1_write),                              //                                          .write
		.btn_s1_readdata                                 (mm_interconnect_0_btn_s1_readdata),                           //                                          .readdata
		.btn_s1_writedata                                (mm_interconnect_0_btn_s1_writedata),                          //                                          .writedata
		.btn_s1_chipselect                               (mm_interconnect_0_btn_s1_chipselect),                         //                                          .chipselect
		.cpu_nios_led3_debug_mem_slave_address           (mm_interconnect_0_cpu_nios_led3_debug_mem_slave_address),     //             cpu_nios_led3_debug_mem_slave.address
		.cpu_nios_led3_debug_mem_slave_write             (mm_interconnect_0_cpu_nios_led3_debug_mem_slave_write),       //                                          .write
		.cpu_nios_led3_debug_mem_slave_read              (mm_interconnect_0_cpu_nios_led3_debug_mem_slave_read),        //                                          .read
		.cpu_nios_led3_debug_mem_slave_readdata          (mm_interconnect_0_cpu_nios_led3_debug_mem_slave_readdata),    //                                          .readdata
		.cpu_nios_led3_debug_mem_slave_writedata         (mm_interconnect_0_cpu_nios_led3_debug_mem_slave_writedata),   //                                          .writedata
		.cpu_nios_led3_debug_mem_slave_byteenable        (mm_interconnect_0_cpu_nios_led3_debug_mem_slave_byteenable),  //                                          .byteenable
		.cpu_nios_led3_debug_mem_slave_waitrequest       (mm_interconnect_0_cpu_nios_led3_debug_mem_slave_waitrequest), //                                          .waitrequest
		.cpu_nios_led3_debug_mem_slave_debugaccess       (mm_interconnect_0_cpu_nios_led3_debug_mem_slave_debugaccess), //                                          .debugaccess
		.jtag_uart_avalon_jtag_slave_address             (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),       //               jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write               (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),         //                                          .write
		.jtag_uart_avalon_jtag_slave_read                (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),          //                                          .read
		.jtag_uart_avalon_jtag_slave_readdata            (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),      //                                          .readdata
		.jtag_uart_avalon_jtag_slave_writedata           (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),     //                                          .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest         (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest),   //                                          .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect          (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),    //                                          .chipselect
		.ledr_s1_address                                 (mm_interconnect_0_ledr_s1_address),                           //                                   ledr_s1.address
		.ledr_s1_write                                   (mm_interconnect_0_ledr_s1_write),                             //                                          .write
		.ledr_s1_readdata                                (mm_interconnect_0_ledr_s1_readdata),                          //                                          .readdata
		.ledr_s1_writedata                               (mm_interconnect_0_ledr_s1_writedata),                         //                                          .writedata
		.ledr_s1_chipselect                              (mm_interconnect_0_ledr_s1_chipselect),                        //                                          .chipselect
		.RAM_s1_address                                  (mm_interconnect_0_ram_s1_address),                            //                                    RAM_s1.address
		.RAM_s1_write                                    (mm_interconnect_0_ram_s1_write),                              //                                          .write
		.RAM_s1_readdata                                 (mm_interconnect_0_ram_s1_readdata),                           //                                          .readdata
		.RAM_s1_writedata                                (mm_interconnect_0_ram_s1_writedata),                          //                                          .writedata
		.RAM_s1_byteenable                               (mm_interconnect_0_ram_s1_byteenable),                         //                                          .byteenable
		.RAM_s1_chipselect                               (mm_interconnect_0_ram_s1_chipselect),                         //                                          .chipselect
		.RAM_s1_clken                                    (mm_interconnect_0_ram_s1_clken),                              //                                          .clken
		.sseg_s1_address                                 (mm_interconnect_0_sseg_s1_address),                           //                                   sseg_s1.address
		.sseg_s1_write                                   (mm_interconnect_0_sseg_s1_write),                             //                                          .write
		.sseg_s1_readdata                                (mm_interconnect_0_sseg_s1_readdata),                          //                                          .readdata
		.sseg_s1_writedata                               (mm_interconnect_0_sseg_s1_writedata),                         //                                          .writedata
		.sseg_s1_chipselect                              (mm_interconnect_0_sseg_s1_chipselect),                        //                                          .chipselect
		.switch_s1_address                               (mm_interconnect_0_switch_s1_address),                         //                                 switch_s1.address
		.switch_s1_readdata                              (mm_interconnect_0_switch_s1_readdata),                        //                                          .readdata
		.sys_timer_s1_address                            (mm_interconnect_0_sys_timer_s1_address),                      //                              sys_timer_s1.address
		.sys_timer_s1_write                              (mm_interconnect_0_sys_timer_s1_write),                        //                                          .write
		.sys_timer_s1_readdata                           (mm_interconnect_0_sys_timer_s1_readdata),                     //                                          .readdata
		.sys_timer_s1_writedata                          (mm_interconnect_0_sys_timer_s1_writedata),                    //                                          .writedata
		.sys_timer_s1_chipselect                         (mm_interconnect_0_sys_timer_s1_chipselect),                   //                                          .chipselect
		.usr_timer_s1_address                            (mm_interconnect_0_usr_timer_s1_address),                      //                              usr_timer_s1.address
		.usr_timer_s1_write                              (mm_interconnect_0_usr_timer_s1_write),                        //                                          .write
		.usr_timer_s1_readdata                           (mm_interconnect_0_usr_timer_s1_readdata),                     //                                          .readdata
		.usr_timer_s1_writedata                          (mm_interconnect_0_usr_timer_s1_writedata),                    //                                          .writedata
		.usr_timer_s1_chipselect                         (mm_interconnect_0_usr_timer_s1_chipselect)                    //                                          .chipselect
	);

	nios_led3_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),       // receiver3.irq
		.sender_irq    (cpu_nios_led3_irq_irq)           //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
